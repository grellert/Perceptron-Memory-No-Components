rom_1_port_v2_inst : rom_1_port_v2 PORT MAP (
		address	 => address_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
