rom_fixedpoint_2048_inst : rom_fixedpoint_2048 PORT MAP (
		address	 => address_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
