rom_fixedpoint_inst : rom_fixedpoint PORT MAP (
		address	 => address_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
